
-- ZX Spectrum Next Hardware Sprites
-- Copyright 2020 Alvin Albrecht
--
-- Sprites v1
-- Theorical Model - Victor Trucco
-- VHDL - Fabio Belavenuto
--
-- Sprites v2
-- Rewritten and enhanced - Alvin Albrecht
-- Ideas - Spectrum Next Team, David Burton, Peter Ped Helcmanovsky
--
-- This file is part of the ZX Spectrum Next Project
-- <https://gitlab.com/SpectrumNext/ZX_Spectrum_Next_FPGA/tree/master/cores>
--
-- The ZX Spectrum Next FPGA source code is free software: you can 
-- redistribute it and/or modify it under the terms of the GNU General 
-- Public License as published by the Free Software Foundation, either 
-- version 3 of the License, or (at your option) any later version.
--
-- The ZX Spectrum Next FPGA source code is distributed in the hope 
-- that it will be useful, but WITHOUT ANY WARRANTY; without even the 
-- implied warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR 
-- PURPOSE.  See the GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with the ZX Spectrum Next FPGA source code.  If not, see 
-- <https://www.gnu.org/licenses/>.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity sprites is
   port (
   
      clock_master_i    : in  std_logic;
      clock_master_180o_i  : in  std_logic;
      clock_pixel_i     : in  std_logic;
      reset_i           : in  std_logic;
      zero_on_top_i     : in  std_logic;
      border_clip_en_i  : in std_logic;
      over_border_i     : in  std_logic;
      hcounter_i        : in  unsigned( 8 downto 0);
      vcounter_i        : in  unsigned( 8 downto 0);
      transp_colour_i   : in  std_logic_vector( 7 downto 0);
      
      -- CPU
      
      port57_w_en_s  : in  std_logic;
      port5B_w_en_s  : in  std_logic;
      port303b_r_en_s: in  std_logic;
      port303b_w_en_s: in  std_logic;
      cpu_d_i        : in  std_logic_vector( 7 downto 0);
      cpu_d_o        : out std_logic_vector( 7 downto 0);
      
      -- NEXTREG MIRROR
      
      mirror_tie_i   : in  std_logic;                       -- 1 = nextreg 0x34 and io port 0x303B tied together
      mirror_we_i    : in  std_logic;
      mirror_index_i : in  std_logic_vector(2 downto 0);    -- attributes 0-4, sprite number if 7
      mirror_data_i  : in  std_logic_vector(7 downto 0);
      mirror_inc_i   : in  std_logic;                       -- one to increment sprite number
      mirror_num_o   : out std_logic_vector(6 downto 0);    -- currently selected sprite number
      
      -- Out
      
      rgb_o          : out std_logic_vector(7 downto 0);
      pixel_en_o     : out std_logic;
      
      -- clip window
      
      clip_x1_i      : in unsigned(7 downto 0);
      clip_x2_i      : in unsigned(7 downto 0);
      clip_y1_i      : in unsigned(7 downto 0);
      clip_y2_i      : in unsigned(7 downto 0)
      
   );
end entity;

architecture rtl of sprites is

   -- the implementation is not fully parameterized primarily because the memories were generated by coregen
   
   constant SPRITE_SIZE_BITS     : integer := 4;  -- sprites are 16x16 pixels
   constant SPRITE_SIZE          : integer := (2 ** SPRITE_SIZE_BITS);
   
-- constant TOTAL_SPRITES_BITS   : integer := 6;  -- 64 sprites total
   constant TOTAL_SPRITES_BITS   : integer := 7;  -- 128 sprites total
   constant TOTAL_SPRITES        : integer := (2 ** TOTAL_SPRITES_BITS);
   
   constant TOTAL_PATTERN_BITS   : integer := 6;  -- 64 different sprite patterns
   constant TOTAL_PATTERNS       : integer := (2 ** TOTAL_PATTERN_BITS);

   -- coregen

   component sdpram_128_8 is
   PORT (

      DPRA  : IN  STD_LOGIC_VECTOR(7-1 downto 0) := (OTHERS => '0');
      CLK   : IN STD_LOGIC;
      WE    : IN  STD_LOGIC;
      DPO   : OUT STD_LOGIC_VECTOR(8-1 downto 0);
      A     : IN  STD_LOGIC_VECTOR(7-1-(4*0*boolean'pos(7>4)) downto 0)
            := (OTHERS => '0');
      D     : IN  STD_LOGIC_VECTOR(8-1 downto 0) := (OTHERS => '0')

   );
   end component;

   component spram_320_9 is
   PORT (

      CLK   : IN STD_LOGIC;
      WE    : IN  STD_LOGIC;
      SPO   : OUT STD_LOGIC_VECTOR(9-1 downto 0);
      A     : IN  STD_LOGIC_VECTOR(9-1-(4*0*boolean'pos(9>4)) downto 0)
            := (OTHERS => '0');
      D     : IN  STD_LOGIC_VECTOR(9-1 downto 0) := (OTHERS => '0')

   );
   end component;

   component sdpbram_16k_8 is
   PORT (
      --Port A
      WEA   : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      ADDRA : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
      DINA  : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      CLKA  : IN STD_LOGIC;
      --Port B
      ENB   : IN STD_LOGIC;  --opt port
      ADDRB : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
      DOUTB : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
      CLKB  : IN STD_LOGIC

   );
   end component;

   -- memory wiring
   
   signal attr_a           : std_logic_vector((TOTAL_SPRITES_BITS-1) downto 0);
   signal attr_id          : std_logic_vector(2 downto 0);
   signal attr_data        : std_logic_vector(7 downto 0);
   signal attr0_we         : std_logic;
   signal attr1_we         : std_logic;
   signal attr2_we         : std_logic;
   signal attr3_we         : std_logic;
   signal attr4_we         : std_logic;
   signal spr_attr_a       : std_logic_vector((TOTAL_SPRITES_BITS-1) downto 0);
   signal sprite_attr_0       : std_logic_vector(7 downto 0);
   signal sprite_attr_1       : std_logic_vector(7 downto 0);
   signal sprite_attr_2    : std_logic_vector(7 downto 0);
   signal sprite_attr_3 : std_logic_vector(7 downto 0);
   signal sprite_attr_4    : std_logic_vector(7 downto 0);
   
   signal l0_we            : std_logic;
   signal l0_a             : std_logic_vector(8 downto 0);
   signal l0_d             : std_logic_vector(8 downto 0);
   signal l0_spo           : std_logic_vector(8 downto 0);
   signal l1_we            : std_logic;
   signal l1_a             : std_logic_vector(8 downto 0);
   signal l1_d             : std_logic_vector(8 downto 0);
   signal l1_spo           : std_logic_vector(8 downto 0);
   signal line_buf_sel     : std_logic;
   
   signal port5b_w_en_d    : std_logic;
   signal pattern_a        : std_logic_vector((TOTAL_PATTERN_BITS+8-1) downto 0);
   signal pattern_we       : std_logic;
   signal spr_pat_addr     : std_logic_vector((TOTAL_PATTERN_BITS+8-1) downto 0);
   signal spr_pat_re       : std_logic;
   signal spr_pat_data     : std_logic_vector(7 downto 0);

   -- cpu port i/o
   
   signal attr_index       : std_logic_vector((TOTAL_SPRITES_BITS+3-1) downto 0);
   signal pattern_index    : std_logic_vector((TOTAL_PATTERN_BITS+8-1) downto 0);
   
   signal index_inc_attr_by_8 : std_logic;
   signal index_inc_in_s      : std_logic_vector((TOTAL_PATTERN_BITS+8-1) downto 0);  -- assumes pattern_index larger than attr_index
   signal index_inc_out_s     : std_logic_vector((TOTAL_PATTERN_BITS+8-1) downto 0);  -- assumes pattern_index larger than attr_index
   
   signal attr_num_change     : std_logic;
   
   signal io_port_access   : std_logic;
   signal io_port_access_d : std_logic;
   signal io_port_re       : std_logic;
   signal cpu_request      : std_logic;
   signal cpu_served       : std_logic;
   signal cpu_sprite_q     : std_logic_vector(TOTAL_SPRITES_BITS-1 downto 0);
   signal cpu_index_q      : std_logic_vector(2 downto 0);
   signal cpu_data_q       : std_logic_vector(7 downto 0);
   
   signal status_reg_s     : std_logic_vector(7 downto 0);
   signal status_reg_read  : std_logic_vector(7 downto 0);
   signal sprites_overtime : std_logic;
   
   -- mirror

   signal mirror_sprite_q  : std_logic_vector(7 downto 0);
   signal mirror_served    : std_logic;
   signal mirror_num_change   : std_logic;
   
   -- load sprite line

   signal line_reset_s     : std_logic;
   signal line_reset_re    : std_logic_vector(1 downto 0);
   signal spr_cur_vcount   : std_logic_vector(8 downto 0);

   signal anchor_rel_type  : std_logic;
   signal anchor_h         : std_logic;
   signal anchor_vis       : std_logic;
   signal anchor_x         : std_logic_vector(8 downto 0);
   signal anchor_y         : std_logic_vector(8 downto 0);
   signal anchor_pattern   : std_logic_vector(6 downto 0);
   signal anchor_paloff    : std_logic_vector(3 downto 0);
   signal anchor_rotate    : std_logic;
   signal anchor_xmirror   : std_logic;
   signal anchor_ymirror   : std_logic;
   signal anchor_xscale    : std_logic_vector(1 downto 0);
   signal anchor_yscale    : std_logic_vector(1 downto 0);

   signal spr_rel_x0       : std_logic_vector(7 downto 0);
   signal spr_rel_y0       : std_logic_vector(7 downto 0);
   signal spr_rel_x1       : std_logic_vector(7 downto 0);
   signal spr_rel_y1       : std_logic_vector(7 downto 0);
   signal spr_rel_x2       : std_logic_vector(8 downto 0);
   signal spr_rel_y2       : std_logic_vector(8 downto 0);
   signal spr_rel_x3       : std_logic_vector(8 downto 0);
   signal spr_rel_y3       : std_logic_vector(8 downto 0);
   
   signal spr_rel_paloff   : std_logic_vector(3 downto 0);
   signal spr_rel_xm       : std_logic;
   signal spr_rel_ym       : std_logic;
   
   signal spr_rel_attr_0   : std_logic_vector(7 downto 0);
   signal spr_rel_attr_1   : std_logic_vector(7 downto 0);
   signal spr_rel_attr_2   : std_logic_vector(7 downto 0);
   signal spr_rel_attr_3   : std_logic_vector(7 downto 0);
   signal spr_rel_attr_4   : std_logic_vector(7 downto 0);
   
   signal spr_cur_attr_0   : std_logic_vector(7 downto 0);
   signal spr_cur_attr_1   : std_logic_vector(7 downto 0);
   signal spr_cur_attr_2   : std_logic_vector(7 downto 0);
   signal spr_cur_attr_3   : std_logic_vector(7 downto 0);
   signal spr_cur_attr_4   : std_logic_vector(7 downto 0);

   signal spr_cur_x        : std_logic_vector(8 downto 0);
   signal spr_cur_y        : std_logic_vector(8 downto 0);
   
   signal spr_relative     : std_logic;
   signal spr_cur_h        : std_logic;
   signal spr_cur_n6       : std_logic;
   signal spr_rel_pattern  : std_logic_vector(6 downto 0);  -- N5:N0,N6
   
   signal spr_y8           : std_logic;
   signal spr_y_offset     : std_logic_vector(8 downto 0);
   signal spr_y_offset_raw : std_logic_vector(8 downto 0);
   signal spr_y_index      : std_logic_vector((SPRITE_SIZE_BITS-1) downto 0);
   signal spr_x_mirr_eff   : std_logic;
   signal spr_x_index      : std_logic_vector((SPRITE_SIZE_BITS-1) downto 0);
   
   signal spr_pattern_addr_start : std_logic_vector((TOTAL_PATTERN_BITS+8-1) downto 0);
   signal spr_pattern_addr_delta : std_logic_vector((TOTAL_PATTERN_BITS+8-1) downto 0);
   
   signal spr_cur_hcount_valid   : std_logic;
   signal spr_cur_notime_mask    : std_logic_vector(4 downto 0);
   signal spr_cur_notime         : std_logic;
   
   signal spr_cur_index          : std_logic_vector((TOTAL_SPRITES_BITS-1) downto 0);
   signal spr_cur_index_is_zero  : std_logic;
   signal spr_width_count        : std_logic_vector((SPRITE_SIZE_BITS-1+1+3) downto 0);
   signal spr_width_count_next   : std_logic_vector((SPRITE_SIZE_BITS-1+1+3) downto 0);
   signal spr_width_count_delta  : std_logic_vector(3 downto 0);
   signal spr_cur_hcount         : std_logic_vector(8 downto 0);
   signal spr_cur_paloff         : std_logic_vector(3 downto 0);
   signal spr_cur_visible        : std_logic;
   signal spr_cur_yoff           : std_logic_vector((8-SPRITE_SIZE_BITS) downto 0);
   signal spr_cur_x_wrap         : std_logic_vector(4 downto 0);
   signal spr_cur_4bit           : std_logic_vector(1 downto 0);
   signal spr_cur_draw_it        : std_logic;
   
   signal spr_cur_pattern_addr   : std_logic_vector((TOTAL_PATTERN_BITS+8-1) downto 0);
   signal spr_cur_pattern_delta  : std_logic_vector((TOTAL_PATTERN_BITS+8-1) downto 0);

   type   state_t          is (S_IDLE, S_START, S_QUALIFY, S_PROCESS);
   signal state_s          : state_t;
   signal state_next_s     : state_t;
   
   signal spr_line_addr_s  : std_logic_vector(8 downto 0);
   signal spr_line_data_s  : std_logic_vector(8 downto 0);
   signal spr_nibble_data  : std_logic_vector(3 downto 0);
   signal spr_line_we      : std_logic;
   signal spr_line_we_s    : std_logic;
   signal spr_line_data_o  : std_logic_vector(8 downto 0);

   -- video line generation
   
   signal hcounter_i_valid : std_logic;
   signal vcounter_i_valid : std_logic;

   signal x_s_v            : unsigned(8 downto 0);
   signal x_e_v            : unsigned(8 downto 0);
   signal y_s_v            : unsigned(8 downto 0);
   signal y_e_v            : unsigned(8 downto 0);
   
   signal over_border_s    : std_logic;

   signal video_line_we_s     : std_logic;
   signal video_line_addr_s   : std_logic_vector(8 downto 0);
   signal video_line_data_s   : std_logic_vector(8 downto 0);
   signal video_line_rgb_s    : std_logic_vector(8 downto 0);
   signal video_line_rgb_load : std_logic_vector(8 downto 0);
   
   signal video_line_re       : std_logic;
   signal video_line_fe       : std_logic;
   signal video_line_flag     : std_logic;

begin

   ----------------------------
   -- SPRITE ATTRIBUTE MEMORIES
   ----------------------------

   -- simple dual port ram (sync write, async read)
   -- X position (bits 7:0)
   
--   attr0 : sdpram_128_8
--   port map (
--      DPRA => spr_attr_a,
--      CLK  => clock_master_180o_i,
--      WE   => attr0_we,
--      DPO  => sprite_attr_0,
--      A    => attr_a,
--      D    => attr_data
--   );

 attr0 : entity work.sdpram
 generic map (
    addr_width_g => TOTAL_SPRITES_BITS,
    data_width_g => 8
 )
 port map (
    clk_a_i  => clock_master_180o_i,
    we_a_i   => attr0_we,
    addr_a_i => attr_a,
    data_a_i => attr_data,
    --
    addr_b_i => spr_attr_a,
    data_b_o => sprite_attr_0
 );

   -- simple dual port ram (sync write, async read)
   -- Y position (bits 7:0)
   
--   attr1 : sdpram_128_8
--   port map (
--      DPRA => spr_attr_a,
--      CLK  => clock_master_180o_i,
--      WE   => attr1_we,
--      DPO  => sprite_attr_1,
--      A    => attr_a,
--      D    => attr_data
--   );

 attr1 : entity work.sdpram
 generic map (
    addr_width_g => TOTAL_SPRITES_BITS,
    data_width_g => 8
 )
 port map (
    clk_a_i  => clock_master_180o_i,
    we_a_i   => attr1_we,
    addr_a_i => attr_a,
    data_a_i => attr_data,
    --
    addr_b_i => spr_attr_a,
    data_b_o => sprite_attr_1
 );

   -- simple dual port ram (sync write, async read)
   -- bits 7-4 is palette offset, bit 3 is X mirror, bit 2 is Y mirror, bit 1 is the rotate flag and bit 0 is X MSB
   
--   attr2 : sdpram_128_8
--   port map (
--      DPRA => spr_attr_a,
--      CLK  => clock_master_180o_i,
--      WE   => attr2_we,
--      DPO  => sprite_attr_2,
--      A    => attr_a,
--      D    => attr_data
--   );

 attr2 : entity work.sdpram
 generic map (
    addr_width_g => TOTAL_SPRITES_BITS,
    data_width_g => 8
 )
 port map (
    clk_a_i  => clock_master_180o_i,
    we_a_i   => attr2_we,
    addr_a_i => attr_a,
    data_a_i => attr_data,
    --
    addr_b_i => spr_attr_a,
    data_b_o => sprite_attr_2
 );

   -- simple dual port ram (sync write, async read)
   -- bit 7 is the visible flag, bit 6 set if fifth attr byte follows, bits 5-0 is Name (pattern index, 0-63)
   
--   attr3 : sdpram_128_8
--   port map (
--      DPRA => spr_attr_a,
--      CLK  => clock_master_180o_i,
--      WE   => attr3_we,
--      DPO  => sprite_attr_3,
--      A    => attr_a,
--      D    => attr_data
--   );

 attr3 : entity work.sdpram
 generic map (
    addr_width_g => TOTAL_SPRITES_BITS,
    data_width_g => 8
 )
 port map (
    clk_a_i  => clock_master_180o_i,
    we_a_i   => attr3_we,
    addr_a_i => attr_a,
    data_a_i => attr_data,
    --
    addr_b_i => spr_attr_a,
    data_b_o => sprite_attr_3
 );

   -- simple dual port ram (sync write, async read)
   -- bit 7 set for 4-bit patterns, bit 6 is Name(6), bit 5 is reserved at 0, bits(4:3) XX scale, bits(2:1) YY scale, bit 0 is Y MSB

--   attr4 : sdpram_128_8
--   port map (
--      DPRA => spr_attr_a,
--      CLK  => clock_master_180o_i,
--      WE   => attr4_we,
--      DPO  => sprite_attr_4,
--      A    => attr_a,
--      D    => attr_data
--   );

 attr4 : entity work.sdpram
 generic map (
    addr_width_g => TOTAL_SPRITES_BITS,
    data_width_g => 8
 )
 port map (
    clk_a_i  => clock_master_180o_i,
    we_a_i   => attr4_we,
    addr_a_i => attr_a,
    data_a_i => attr_data,
    --
    addr_b_i => spr_attr_a,
    data_b_o => sprite_attr_4
 );

   -----------------------------
   -- VIDEO LINE BUFFER MEMORIES
   -----------------------------

   -- single port ram (sync write, async read)
   
--   linebuf0 : spram_320_9
--   port map (
--      CLK  => clock_master_180o_i,
--      WE   => l0_we,
--      SPO  => l0_spo,
--      A    => l0_a,
--      D    => l0_d
--   );

 linebuf0 : entity work.spram
 generic map (
    addr_width_g => 9,
    data_width_g => 9
 )
 port map (
    clk_i    => clock_master_180o_i,
    we_i     => l0_we,
    addr_i   => l0_a,
    data_i   => l0_d,
    data_o   => l0_spo
 );

   -- single port ram (sync write, async read)
   
--   linebuf1 : spram_320_9
--   port map (
--      CLK  => clock_master_180o_i,
--      WE   => l1_we,
--      SPO  => l1_spo,
--      A    => l1_a,
--      D    => l1_d
--   );

 linebuf1 : entity work.spram
 generic map (
    addr_width_g => 9,
    data_width_g => 9
 )
 port map (
    clk_i    => clock_master_180o_i,
    we_i     => l1_we,
    addr_i   => l1_a,
    data_i   => l1_d,
    data_o   => l1_spo
 );

   -- swap line buffers between sprite and video
   
   line_reset_s <= '1' when hcounter_i = "111111111" else '0';
   
   process (clock_master_i)
   begin
      if rising_edge(clock_master_i) then
         if reset_i = '1' then
            line_reset_re <= "00";
         else
            line_reset_re <= line_reset_re(0) & line_reset_s;
         end if;
      end if;
   end process;
   
   process (clock_master_i)
   begin
      if rising_edge(clock_master_i) then
         if reset_i = '1' then
            line_buf_sel <= '0';
            spr_cur_vcount <= (others => '0');
         elsif line_reset_re = "01" then
            line_buf_sel <= not line_buf_sel;
            spr_cur_vcount <= std_logic_vector(vcounter_i + 1);
         end if;
      end if;
   end process;
   
   l0_we <= video_line_we_s   when line_buf_sel = '0' else spr_line_we_s;
   l0_a  <= video_line_addr_s when line_buf_sel = '0' else spr_line_addr_s;
   l0_d  <= video_line_data_s when line_buf_sel = '0' else spr_line_data_s;
   
   l1_we <= spr_line_we_s     when line_buf_sel = '0' else video_line_we_s;
   l1_a  <= spr_line_addr_s   when line_buf_sel = '0' else video_line_addr_s;
   l1_d  <= spr_line_data_s   when line_buf_sel = '0' else video_line_data_s;
   
   spr_line_data_o  <= l1_spo when line_buf_sel = '0' else l0_spo;
   video_line_rgb_s <= l0_spo when line_buf_sel = '0' else l1_spo;
   
   -----------------
   -- PATTERN MEMORY
   -----------------
   
   -- simple dual port ram (sync write, sync read zero delay)
   
--   pattern : sdpbram_16k_8
--   port map (
--      WEA        => pattern_we,
--      ADDRA      => pattern_a,
--      DINA       => cpu_data_q,
--      CLKA       => clock_master_180o_i,
--      --
--      ENB        => '1', 
--      ADDRB      => spr_pat_addr,
--      DOUTB      => spr_pat_data,
--      CLKB       => clock_master_i
--   );

 pattern: entity work.dpram
 generic map (
    addr_width_g => (TOTAL_SPRITES_BITS+7),
    data_width_g => 8
 )
 port map (
    clk_a_i  => clock_master_180o_i,
    we_i     => pattern_we,
    addr_a_i => pattern_a,
    data_a_i => cpu_data_q,
    --
    clk_b_i  => clock_master_i,
    addr_b_i => spr_pat_addr,
    data_b_o => spr_pat_data
 );

   -----------------
   -- NEXTREG MIRROR
   -----------------
   
   process (clock_master_i)
   begin
      if rising_edge(clock_master_i) then
         mirror_num_change <= '0';
         if reset_i = '1' then
            mirror_sprite_q <= (others => '0');
         elsif mirror_we_i = '1' and mirror_index_i = "111" then
            mirror_sprite_q <= mirror_data_i;
            mirror_num_change <= '1';
         elsif mirror_inc_i = '1' then
            mirror_sprite_q(TOTAL_SPRITES_BITS-1 downto 0) <= mirror_sprite_q(TOTAL_SPRITES_BITS-1 downto 0) + 1;
            mirror_sprite_q(7) <= pattern_index(7);
            mirror_num_change <= '1';
         elsif attr_num_change = '1' and mirror_tie_i = '1' then
            mirror_sprite_q(TOTAL_SPRITES_BITS-1 downto 0) <= attr_index((TOTAL_SPRITES_BITS+3-1) downto 3);
            mirror_sprite_q(7) <= pattern_index(7);   -- wear helmet
         end if;
      end if;
   end process;

   mirror_num_o <= mirror_sprite_q(TOTAL_SPRITES_BITS-1 downto 0);

   ----------------------
   -- CPU SPRITE PORT I/O
   ----------------------
   
   -- rising edge detection
   
   io_port_access <= '1' when port57_w_en_s = '1' or port5B_w_en_s = '1' or port303b_r_en_s = '1' or port303b_w_en_s = '1' else '0';
   
   process (clock_master_i)
   begin
      if rising_edge(clock_master_i) then
         if reset_i = '1' then
            io_port_access_d <= '0';
         else
            io_port_access_d <= io_port_access;
         end if;
      end if;
   end process;
   
   io_port_re <= io_port_access and not io_port_access_d;

   -- cpu ports 0x57, 0x5b, 0x303b
   
   index_inc_attr_by_8 <= '1' when attr_index(2) = '1' or (attr_index(2 downto 0) = "011" and cpu_d_i(6) = '0') else '0';

   index_inc_in_s <= ("0000" & attr_index) when port57_w_en_s = '1' and index_inc_attr_by_8 = '0' else
                     ("0000000" & attr_index((TOTAL_SPRITES_BITS+3-1) downto 3)) when port57_w_en_s = '1' and index_inc_attr_by_8 = '1' else
                     pattern_index;

   index_inc_out_s <= index_inc_in_s + 1;
   
   process (clock_master_i)
   begin
      if rising_edge(clock_master_i) then
         attr_num_change <= '0';
         if reset_i = '1' then
            attr_index <= (others => '0');
         elsif mirror_num_change = '1' and mirror_tie_i = '1' then
            attr_index <= mirror_sprite_q(TOTAL_SPRITES_BITS-1 downto 0) & "000";
         elsif port303b_w_en_s = '1' and io_port_re = '1' then
            attr_index <= cpu_d_i(TOTAL_SPRITES_BITS-1 downto 0) & "000";
            attr_num_change <= '1';
         elsif port57_w_en_s = '1' and io_port_re = '1' then
            if index_inc_attr_by_8 = '0' then
               attr_index <= index_inc_out_s((TOTAL_SPRITES_BITS+3-1) downto 0);
            else
               attr_index <= index_inc_out_s((TOTAL_SPRITES_BITS-1) downto 0) & "000";
               attr_num_change <= '1';
            end if;
         end if;
      end if;
   end process;

   process (clock_master_i)
   begin
      if rising_edge(clock_master_i) then
         if reset_i = '1' then
            cpu_sprite_q <= (others => '0');
            cpu_index_q <= (others => '0');
         elsif port57_w_en_s = '1' and io_port_re = '1' then
            cpu_sprite_q <= attr_index((TOTAL_SPRITES_BITS+3-1) downto 3);
            cpu_index_q <= attr_index(2 downto 0);
         end if;
      end if;
   end process;
   
   process (clock_master_i)
   begin
      if rising_edge(clock_master_i) then
         if io_port_re = '1' then
            cpu_data_q <= cpu_d_i;
         end if;
      end if;
   end process;
   
   process (clock_master_i)
   begin
      if rising_edge(clock_master_i) then
         if reset_i = '1' then
            cpu_request <= '0';
         elsif port57_w_en_s = '1' and io_port_re = '1' then
            cpu_request <= '1';
         elsif cpu_served = '1' then
            cpu_request <= '0';
         end if;
      end if;
   end process;

   mirror_served <= '1' when mirror_we_i = '1' and mirror_index_i <= "100" else '0';
   cpu_served <= '1' when mirror_served = '0' and cpu_request = '1' else '0';

   attr_a    <= cpu_sprite_q when mirror_served = '0' else mirror_sprite_q(TOTAL_SPRITES_BITS-1 downto 0);
   attr_id   <= cpu_index_q when mirror_served = '0' else mirror_index_i;
   attr_data <= cpu_data_q when mirror_served = '0' else mirror_data_i;
   
   attr0_we <= '1' when (cpu_served = '1' or mirror_served = '1') and attr_id = "000" else '0';
   attr1_we <= '1' when (cpu_served = '1' or mirror_served = '1') and attr_id = "001" else '0';
   attr2_we <= '1' when (cpu_served = '1' or mirror_served = '1') and attr_id = "010" else '0';
   attr3_we <= '1' when (cpu_served = '1' or mirror_served = '1') and attr_id = "011" else '0';
   attr4_we <= '1' when (cpu_served = '1' or mirror_served = '1') and attr_id = "100" else '0';
   
   process (clock_master_i)
   begin
      if rising_edge(clock_master_i) then
         if reset_i = '1' then
            port5b_w_en_d <= '0';
         else
            port5b_w_en_d <= port5b_w_en_s and io_port_re;
         end if;
      end if;
   end process;
   
   process (clock_master_i)
   begin
      if rising_edge(clock_master_i) then
         if reset_i = '1' then
            pattern_index <= (others => '0');
         elsif mirror_num_change = '1' and mirror_tie_i = '1' then
            pattern_index <= mirror_sprite_q(TOTAL_PATTERN_BITS-1 downto 0) & mirror_sprite_q(7) & "0000000";
         elsif port303b_w_en_s = '1' and io_port_re = '1' then
            pattern_index <= cpu_d_i(TOTAL_PATTERN_BITS-1 downto 0) & cpu_d_i(7) & "0000000";
         elsif port5b_w_en_d = '1' then
            pattern_index <= index_inc_out_s;
         end if;
      end if;
   end process;

   pattern_a <= pattern_index;
   pattern_we <= '1' when port5b_w_en_d = '1' else '0';
   
   -- cpu port 0x303b read

   cpu_d_o <= status_reg_read;
   
   -------------------
   -- LOAD SPRITE LINE
   -------------------
   
   -- maybe there is a better way to do this
   
   spr_relative <= '1' when sprite_attr_3(6) = '1' and sprite_attr_4(7 downto 6) = "01" else '0';

   -- sort out relative sprite characteristics
   
   spr_rel_x0 <= sprite_attr_0 when anchor_rotate = '0' else sprite_attr_1;
   spr_rel_y0 <= sprite_attr_1 when anchor_rotate = '0' else sprite_attr_0;
   spr_rel_x1 <= spr_rel_x0 when (anchor_rotate xor anchor_xmirror) = '0' else (not(spr_rel_x0) + 1);
   spr_rel_y1 <= spr_rel_y0 when anchor_ymirror = '0' else (not(spr_rel_y0) + 1);
   spr_rel_x2 <= (spr_rel_x1(7) & spr_rel_x1)      when anchor_xscale = "00" else
                 (spr_rel_x1 & '0')                when anchor_xscale = "01" else
                 (spr_rel_x1(6 downto 0) & "00")   when anchor_xscale = "10" else
                 (spr_rel_x1(5 downto 0) & "000");
   spr_rel_y2 <= (spr_rel_y1(7) & spr_rel_y1)      when anchor_yscale = "00" else
                 (spr_rel_y1 & '0')                when anchor_yscale = "01" else
                 (spr_rel_y1(6 downto 0) & "00")   when anchor_yscale = "10" else
                 (spr_rel_y1(5 downto 0) & "000");
   spr_rel_x3 <= anchor_x + spr_rel_x2;
   spr_rel_y3 <= anchor_y + spr_rel_y2;
   
   spr_rel_paloff <= sprite_attr_2(7 downto 4) when sprite_attr_2(0) = '0' else (anchor_paloff + sprite_attr_2(7 downto 4));
   
   spr_rel_xm <= sprite_attr_2(3) when anchor_rotate = '0' else sprite_attr_2(2) xor sprite_attr_2(1);
   spr_rel_ym <= sprite_attr_2(2) when anchor_rotate = '0' else sprite_attr_2(3) xor sprite_attr_2(1);

   spr_rel_attr_0 <= spr_rel_x3(7 downto 0);
   spr_rel_attr_1 <= spr_rel_y3(7 downto 0);
   spr_rel_attr_2 <= (spr_rel_paloff & sprite_attr_2(3 downto 1) & spr_rel_x3(8)) when anchor_rel_type = '0' else
                     (spr_rel_paloff & (anchor_xmirror xor spr_rel_xm) & (anchor_ymirror xor spr_rel_ym) & (anchor_rotate xor sprite_attr_2(1)) & spr_rel_x3(8));
   spr_rel_attr_3 <= (anchor_vis and sprite_attr_3(7)) & '1' & sprite_attr_3(5 downto 0);
   spr_rel_attr_4 <= (anchor_h & sprite_attr_4(5) & '0' & sprite_attr_4(4 downto 1) & spr_rel_y3(8)) when anchor_rel_type = '0' else
                     (anchor_h & sprite_attr_4(5) & '0' & anchor_xscale & anchor_yscale & spr_rel_y3(8));

   spr_cur_attr_0 <= sprite_attr_0 when spr_relative = '0' else spr_rel_attr_0;
   spr_cur_attr_1 <= sprite_attr_1 when spr_relative = '0' else spr_rel_attr_1;
   spr_cur_attr_2 <= sprite_attr_2 when spr_relative = '0' else spr_rel_attr_2;
   spr_cur_attr_3 <= sprite_attr_3 when spr_relative = '0' else spr_rel_attr_3;
   spr_cur_attr_4 <= sprite_attr_4 when spr_relative = '0' else spr_rel_attr_4;
   
   -- sprite processing

   spr_y8 <= '0' when sprite_attr_3(6) = '0' else spr_cur_attr_4(0);
   spr_cur_y <= spr_y8 & spr_cur_attr_1;
   
   spr_cur_x <= spr_cur_attr_2(0) & spr_cur_attr_0;
   
   spr_cur_h <= spr_cur_attr_4(7) and sprite_attr_3(6);
   spr_cur_n6 <= spr_cur_attr_4(6) and spr_cur_h;
   spr_rel_pattern <= ((sprite_attr_3((TOTAL_PATTERN_BITS-1) downto 0) & spr_cur_n6) + anchor_pattern) when (spr_relative = '1') and (sprite_attr_4(0) = '1') else
                       (sprite_attr_3((TOTAL_PATTERN_BITS-1) downto 0) & spr_cur_n6);
   
   spr_y_offset_raw <= spr_cur_vcount - spr_cur_y;
   spr_y_offset <= spr_y_offset_raw when sprite_attr_3(6) = '0' or spr_cur_attr_4(2 downto 1) = "00" else
                   spr_y_offset_raw(8) & spr_y_offset_raw(8 downto 1) when spr_cur_attr_4(2 downto 1) = "01" else
                   spr_y_offset_raw(8) & spr_y_offset_raw(8) & spr_y_offset_raw(8 downto 2) when spr_cur_attr_4(2 downto 1) = "10" else
                   spr_y_offset_raw(8) & spr_y_offset_raw(8) & spr_y_offset_raw(8) & spr_y_offset_raw(8 downto 3);
   spr_y_index <= spr_y_offset((SPRITE_SIZE_BITS-1) downto 0) when spr_cur_attr_2(2) = '0' else not(spr_y_offset((SPRITE_SIZE_BITS-1) downto 0));   -- complement for y mirror
   
   spr_x_mirr_eff <= spr_cur_attr_2(3) xor spr_cur_attr_2(1);  -- rotation inverts x mirror
   spr_x_index <= std_logic_vector(to_unsigned(0,spr_x_index'length)) when spr_x_mirr_eff = '0' else std_logic_vector(to_unsigned(65535,spr_x_index'length));
   
   spr_pattern_addr_start <= (spr_rel_pattern(TOTAL_PATTERN_BITS downto 1) & spr_y_index & spr_x_index) when spr_cur_attr_2(1) = '0' else (spr_rel_pattern(TOTAL_PATTERN_BITS downto 1) & spr_x_index & spr_y_index);  -- rotation
   spr_pattern_addr_delta <= "11" & X"FF0" when spr_x_mirr_eff = '1' and spr_cur_attr_2(1) = '1' else  -- x mirror and rotate: -16
                             "11" & X"FFF" when spr_x_mirr_eff = '1' and spr_cur_attr_2(1) = '0' else  -- x mirror and no rotate: -1
                             "00" & X"010" when spr_x_mirr_eff = '0' and spr_cur_attr_2(1) = '1' else  -- no x mirror and rotate: +16
                             "00" & X"001";
   
   spr_cur_hcount_valid <= '1' when spr_cur_hcount < 320 else '0';
   
   spr_cur_notime_mask <= spr_cur_x_wrap(2 downto 0) & "00";
   spr_cur_notime <= '1' when hcounter_i_valid = '1' and hcounter_i(8) = '1' and hcounter_i(5) = '1' and ((std_logic_vector(hcounter_i(4 downto 0)) and spr_cur_notime_mask) = spr_cur_notime_mask) else '0';

   -- state
   
   process (clock_master_i)
   begin
      if rising_edge(clock_master_i) then
         if reset_i = '1' then
            state_s <= S_IDLE;
         elsif line_reset_re = "01" then
            state_s <= S_START;
         else
            state_s <= state_next_s;
         end if;
      end if;
   end process;
   
   -- next state combinatorial
   
   spr_cur_index_is_zero <= '1' when spr_cur_index = 0 else '0';
   spr_cur_draw_it <= '1' when spr_cur_visible = '1' and spr_cur_yoff = 0 else '0';
   
   process (state_s, spr_cur_draw_it, spr_cur_index_is_zero, spr_width_count, spr_cur_hcount_valid, spr_cur_hcount, spr_cur_x_wrap, spr_cur_notime)
   begin
      case state_s is
         when S_START   => state_next_s <= S_QUALIFY;
         when S_QUALIFY => if spr_cur_draw_it = '1' and spr_cur_notime = '1' then
                              state_next_s <= S_IDLE;
                           elsif spr_cur_draw_it = '1' then
                              state_next_s <= S_PROCESS;
                           elsif spr_cur_index_is_zero = '1' then
                              state_next_s <= S_IDLE;
                           else
                              state_next_s <= S_QUALIFY;
                           end if;
         when S_PROCESS => if spr_width_count(SPRITE_SIZE_BITS-1+1+3) = '1' or (spr_cur_hcount_valid = '0' and ((spr_cur_hcount(8 downto 4) and spr_cur_x_wrap) /= spr_cur_x_wrap)) then   -- allow x wrap-around
                              if spr_cur_index_is_zero = '1' then
                                 state_next_s <= S_IDLE;
                              else
                                 state_next_s <= S_QUALIFY;
                              end if;
                           else
                              state_next_s <= S_PROCESS;
                           end if;
         when others    => state_next_s <= S_IDLE;
      end case;
   end process;

   -- state machine variables

   spr_width_count_next <= spr_width_count + spr_width_count_delta;
   
   process (clock_master_180o_i)
   begin
      if rising_edge(clock_master_180o_i) then
         if reset_i = '1' then
            spr_cur_index <= (others => '0');
            spr_cur_hcount <= (others => '0');
            spr_cur_pattern_addr <= (others => '0');
            spr_cur_pattern_delta <= (others => '0');
            spr_width_count <= (others => '0');
            spr_cur_paloff <= (others => '0');
            spr_cur_visible <= '0';
            spr_cur_yoff <= (others => '0');
            spr_cur_x_wrap <= (others => '0');
            spr_cur_4bit <= (others => '0');
            anchor_rel_type <= '0';
            anchor_h <= '0';
            anchor_vis <= '0';
            anchor_x <= (others => '0');
            anchor_y <= (others => '0');
            anchor_pattern <= (others => '0');
            anchor_paloff <= (others => '0');
            anchor_rotate <= '0';
            anchor_xmirror <= '0';
            anchor_ymirror <= '0';
            anchor_xscale <= (others => '0');
            anchor_yscale <= (others => '0');
         elsif state_s = S_START then
            spr_cur_index <= (others => '0');
            anchor_vis <= '0';
         elsif state_s = S_QUALIFY then
            spr_cur_index <= spr_cur_index + 1;
            spr_cur_hcount <= spr_cur_x;
            spr_cur_pattern_addr <= spr_pattern_addr_start;
            spr_cur_pattern_delta <= spr_pattern_addr_delta;
            spr_width_count <= (others => '0');
            if sprite_attr_3(6) = '0' or spr_cur_attr_4(4 downto 3) = "00" then
               spr_width_count_delta <= "1000";
            elsif spr_cur_attr_4(4 downto 3) = "01" then
               spr_width_count_delta <= "0100";
            elsif spr_cur_attr_4(4 downto 3) = "10" then
               spr_width_count_delta <= "0010";
            else
               spr_width_count_delta <= "0001";
            end if;
            spr_cur_paloff <= spr_cur_attr_2(7 downto 4);
            spr_cur_visible <= spr_cur_attr_3(7);
            spr_cur_yoff <= spr_y_offset(8 downto SPRITE_SIZE_BITS);
            if sprite_attr_3(6) = '0' or spr_cur_attr_4(4 downto 3) = "00" then
               spr_cur_x_wrap <= "11111";
            elsif spr_cur_attr_4(4 downto 3) = "01" then
               spr_cur_x_wrap <= "11110";
            elsif spr_cur_attr_4(4 downto 3) = "10" then
               spr_cur_x_wrap <= "11100";
            else
               spr_cur_x_wrap <= "11000";
            end if;
            spr_cur_4bit <= spr_cur_h & spr_rel_pattern(0);
            if spr_relative = '0' then
               anchor_rel_type <= sprite_attr_4(5) and sprite_attr_3(6);
               anchor_h <= sprite_attr_4(7) and sprite_attr_3(6);
               anchor_vis <= sprite_attr_3(7);
               anchor_x <= spr_cur_x;
               anchor_y <= spr_cur_y;
               anchor_pattern <= spr_rel_pattern;
               anchor_paloff <= sprite_attr_2(7 downto 4);
               if sprite_attr_3(6) = '1' and sprite_attr_4(5) = '1' then
                  anchor_rotate <= sprite_attr_2(1);
                  anchor_xmirror <= sprite_attr_2(3);
                  anchor_ymirror <= sprite_attr_2(2);
                  anchor_xscale <= sprite_attr_4(4 downto 3);
                  anchor_yscale <= sprite_attr_4(2 downto 1);
               else
                  anchor_rotate <= '0';
                  anchor_xmirror <= '0';
                  anchor_ymirror <= '0';
                  anchor_xscale <= "00";
                  anchor_yscale <= "00";
               end if;
            end if;
         elsif state_s = S_PROCESS then
            spr_width_count <= spr_width_count_next;
            spr_cur_hcount <= spr_cur_hcount + 1;
            if spr_width_count_next(3) /= spr_width_count(3) then
               spr_cur_pattern_addr <= spr_cur_pattern_addr + spr_cur_pattern_delta;
            end if;
         end if;
      end if;
   end process;

   spr_attr_a <= spr_cur_index;
   spr_pat_addr <= spr_cur_pattern_addr when spr_cur_4bit(1) = '0' else
                   spr_cur_pattern_addr(13 downto 8) & spr_cur_4bit(0) & spr_cur_pattern_addr(7 downto 1);

   spr_line_addr_s <= spr_cur_hcount;

   spr_nibble_data <= spr_pat_data(7 downto 4) when spr_cur_pattern_addr(0) = '0' else spr_pat_data(3 downto 0);
   spr_line_data_s(7 downto 0) <= ((spr_pat_data(7 downto 4) + spr_cur_paloff) & spr_pat_data(3 downto 0)) when spr_cur_4bit(1) = '0' else (spr_cur_paloff & spr_nibble_data(3 downto 0));
   spr_line_data_s(8) <= '1';

   spr_line_we <= '1' when state_s = S_PROCESS and spr_cur_hcount_valid = '1' and ((spr_cur_4bit(1) = '0' and spr_pat_data(7 downto 0) /= transp_colour_i) or (spr_cur_4bit(1) = '1' and spr_nibble_data /= transp_colour_i(3 downto 0))) else '0';
   spr_line_we_s <= '1' when spr_line_we = '1' and (zero_on_top_i = '0' or spr_line_data_o(8) = '0') else '0';

   -- status register
   -- bits(7:2) = 0, bit 1 = max sprites per line, bit 0 = collision 

   process (clock_master_i)
   begin
      if rising_edge(clock_master_i) then
         if reset_i = '1' then
            sprites_overtime <= '0';
         elsif (state_s /= S_IDLE and line_reset_re = "01") or (state_s = S_QUALIFY and spr_cur_notime = '1' and spr_cur_draw_it = '1') then
            sprites_overtime <= '1';
         else
            sprites_overtime <= '0';
         end if;
      end if;
   end process;
   
   process (clock_master_180o_i)
   begin
      if rising_edge(clock_master_180o_i) then
         if (reset_i = '1') then
            status_reg_s <= (others => '0');
            status_reg_read <= (others => '0');
         else
            if port303b_r_en_s = '1' and io_port_re = '1' then
               status_reg_read <= status_reg_s;
               status_reg_s <= (others => '0');
            else
               status_reg_s(1) <= status_reg_s(1) or sprites_overtime;
               status_reg_s(0) <= status_reg_s(0) or (spr_line_data_o(8) and spr_line_we);
            end if;
         end if;
      end if;
   end process;

   -----------------------------
   -- GENERATE VIDEO LINE OUTPUT
   -----------------------------
   
   hcounter_i_valid <= '1' when hcounter_i < 320 else '0';
   vcounter_i_valid <= '1' when vcounter_i(8) = '0' else '0';   -- < 256

   process (clock_pixel_i)
   begin
      if rising_edge(clock_pixel_i) then
         if reset_i = '1' then
            video_line_flag <= '0';
         else
            video_line_flag <= not(video_line_flag);
         end if;
      end if;
   end process;

   -- load video line pixel before clearing
   
   process (clock_pixel_i)
   begin
      if falling_edge(clock_pixel_i) then
         if reset_i = '1' then
            video_line_rgb_load <= (others => '0');
         else
            video_line_rgb_load <= video_line_rgb_s;
            video_line_fe <= video_line_flag;
         end if;
      end if;
   end process;
   
   -- clear video line pixel after loaded
   
   video_line_we_s <= (video_line_fe xor video_line_re) and hcounter_i_valid;
   video_line_addr_s <= std_logic_vector(hcounter_i);
   video_line_data_s <= std_logic_vector(to_unsigned(0,video_line_data_s'length));
   
   -- send video line pixel to display
   
   process (clock_pixel_i)
   begin
      if rising_edge(clock_pixel_i) then
      
         video_line_re <= video_line_flag;

         if over_border_i = '1' then
            if border_clip_en_i = '0' then
               x_s_v <= to_unsigned(0,   9);
               x_e_v <= to_unsigned(319, 9);
               y_s_v <= to_unsigned(0,   9);
               y_e_v <= to_unsigned(255, 9);
            else
               x_s_v <= clip_x1_i & '0';
               x_e_v <= clip_x2_i & '1';
               y_s_v <= '0' & clip_y1_i;
               y_e_v <= '0' & clip_y2_i;
            end if;
         else
            x_s_v <= (('0' & clip_x1_i(7 downto 5)) + 1) & clip_x1_i(4 downto 0);
            x_e_v <= (('0' & clip_x2_i(7 downto 5)) + 1) & clip_x2_i(4 downto 0);
            y_s_v <= (('0' & clip_y1_i(7 downto 5)) + 1) & clip_y1_i(4 downto 0);
            y_e_v <= (('0' & clip_y2_i(7 downto 5)) + 1) & clip_y2_i(4 downto 0);
         end if;
         
         over_border_s <= over_border_i;
      
      end if;
   end process;

   pixel_en_o <= video_line_rgb_load(8) when (vcounter_i >= y_s_v and vcounter_i <= y_e_v and (over_border_s = '1' or vcounter_i < 224) and hcounter_i >= x_s_v and hcounter_i <= x_e_v and hcounter_i_valid = '1' and vcounter_i_valid = '1') else '0';
   rgb_o <= video_line_rgb_load(7 downto 0);

end architecture;
